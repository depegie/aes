module aes_inv_sbox (
    input      [7 : 0] input_byte,
    output reg [7 : 0] output_byte
);
    always_comb begin
        case (input_byte)
    		8'h00: output_byte = 8'h52;
			8'h01: output_byte = 8'h09;
			8'h02: output_byte = 8'h6a;
			8'h03: output_byte = 8'hd5;
			8'h04: output_byte = 8'h30;
			8'h05: output_byte = 8'h36;
			8'h06: output_byte = 8'ha5;
			8'h07: output_byte = 8'h38;
			8'h08: output_byte = 8'hbf;
			8'h09: output_byte = 8'h40;
			8'h0a: output_byte = 8'ha3;
			8'h0b: output_byte = 8'h9e;
			8'h0c: output_byte = 8'h81;
			8'h0d: output_byte = 8'hf3;
			8'h0e: output_byte = 8'hd7;
			8'h0f: output_byte = 8'hfb;
			8'h10: output_byte = 8'h7c;
			8'h11: output_byte = 8'he3;
			8'h12: output_byte = 8'h39;
			8'h13: output_byte = 8'h82;
			8'h14: output_byte = 8'h9b;
			8'h15: output_byte = 8'h2f;
			8'h16: output_byte = 8'hff;
			8'h17: output_byte = 8'h87;
			8'h18: output_byte = 8'h34;
			8'h19: output_byte = 8'h8e;
			8'h1a: output_byte = 8'h43;
			8'h1b: output_byte = 8'h44;
			8'h1c: output_byte = 8'hc4;
			8'h1d: output_byte = 8'hde;
			8'h1e: output_byte = 8'he9;
			8'h1f: output_byte = 8'hcb;
			8'h20: output_byte = 8'h54;
			8'h21: output_byte = 8'h7b;
			8'h22: output_byte = 8'h94;
			8'h23: output_byte = 8'h32;
			8'h24: output_byte = 8'ha6;
			8'h25: output_byte = 8'hc2;
			8'h26: output_byte = 8'h23;
			8'h27: output_byte = 8'h3d;
			8'h28: output_byte = 8'hee;
			8'h29: output_byte = 8'h4c;
			8'h2a: output_byte = 8'h95;
			8'h2b: output_byte = 8'h0b;
			8'h2c: output_byte = 8'h42;
			8'h2d: output_byte = 8'hfa;
			8'h2e: output_byte = 8'hc3;
			8'h2f: output_byte = 8'h4e;
			8'h30: output_byte = 8'h08;
			8'h31: output_byte = 8'h2e;
			8'h32: output_byte = 8'ha1;
			8'h33: output_byte = 8'h66;
			8'h34: output_byte = 8'h28;
			8'h35: output_byte = 8'hd9;
			8'h36: output_byte = 8'h24;
			8'h37: output_byte = 8'hb2;
			8'h38: output_byte = 8'h76;
			8'h39: output_byte = 8'h5b;
			8'h3a: output_byte = 8'ha2;
			8'h3b: output_byte = 8'h49;
			8'h3c: output_byte = 8'h6d;
			8'h3d: output_byte = 8'h8b;
			8'h3e: output_byte = 8'hd1;
			8'h3f: output_byte = 8'h25;
			8'h40: output_byte = 8'h72;
			8'h41: output_byte = 8'hf8;
			8'h42: output_byte = 8'hf6;
			8'h43: output_byte = 8'h64;
			8'h44: output_byte = 8'h86;
			8'h45: output_byte = 8'h68;
			8'h46: output_byte = 8'h98;
			8'h47: output_byte = 8'h16;
			8'h48: output_byte = 8'hd4;
			8'h49: output_byte = 8'ha4;
			8'h4a: output_byte = 8'h5c;
			8'h4b: output_byte = 8'hcc;
			8'h4c: output_byte = 8'h5d;
			8'h4d: output_byte = 8'h65;
			8'h4e: output_byte = 8'hb6;
			8'h4f: output_byte = 8'h92;
			8'h50: output_byte = 8'h6c;
			8'h51: output_byte = 8'h70;
			8'h52: output_byte = 8'h48;
			8'h53: output_byte = 8'h50;
			8'h54: output_byte = 8'hfd;
			8'h55: output_byte = 8'hed;
			8'h56: output_byte = 8'hb9;
			8'h57: output_byte = 8'hda;
			8'h58: output_byte = 8'h5e;
			8'h59: output_byte = 8'h15;
			8'h5a: output_byte = 8'h46;
			8'h5b: output_byte = 8'h57;
			8'h5c: output_byte = 8'ha7;
			8'h5d: output_byte = 8'h8d;
			8'h5e: output_byte = 8'h9d;
			8'h5f: output_byte = 8'h84;
			8'h60: output_byte = 8'h90;
			8'h61: output_byte = 8'hd8;
			8'h62: output_byte = 8'hab;
			8'h63: output_byte = 8'h00;
			8'h64: output_byte = 8'h8c;
			8'h65: output_byte = 8'hbc;
			8'h66: output_byte = 8'hd3;
			8'h67: output_byte = 8'h0a;
			8'h68: output_byte = 8'hf7;
			8'h69: output_byte = 8'he4;
			8'h6a: output_byte = 8'h58;
			8'h6b: output_byte = 8'h05;
			8'h6c: output_byte = 8'hb8;
			8'h6d: output_byte = 8'hb3;
			8'h6e: output_byte = 8'h45;
			8'h6f: output_byte = 8'h06;
			8'h70: output_byte = 8'hd0;
			8'h71: output_byte = 8'h2c;
			8'h72: output_byte = 8'h1e;
			8'h73: output_byte = 8'h8f;
			8'h74: output_byte = 8'hca;
			8'h75: output_byte = 8'h3f;
			8'h76: output_byte = 8'h0f;
			8'h77: output_byte = 8'h02;
			8'h78: output_byte = 8'hc1;
			8'h79: output_byte = 8'haf;
			8'h7a: output_byte = 8'hbd;
			8'h7b: output_byte = 8'h03;
			8'h7c: output_byte = 8'h01;
			8'h7d: output_byte = 8'h13;
			8'h7e: output_byte = 8'h8a;
			8'h7f: output_byte = 8'h6b;
			8'h80: output_byte = 8'h3a;
			8'h81: output_byte = 8'h91;
			8'h82: output_byte = 8'h11;
			8'h83: output_byte = 8'h41;
			8'h84: output_byte = 8'h4f;
			8'h85: output_byte = 8'h67;
			8'h86: output_byte = 8'hdc;
			8'h87: output_byte = 8'hea;
			8'h88: output_byte = 8'h97;
			8'h89: output_byte = 8'hf2;
			8'h8a: output_byte = 8'hcf;
			8'h8b: output_byte = 8'hce;
			8'h8c: output_byte = 8'hf0;
			8'h8d: output_byte = 8'hb4;
			8'h8e: output_byte = 8'he6;
			8'h8f: output_byte = 8'h73;
			8'h90: output_byte = 8'h96;
			8'h91: output_byte = 8'hac;
			8'h92: output_byte = 8'h74;
			8'h93: output_byte = 8'h22;
			8'h94: output_byte = 8'he7;
			8'h95: output_byte = 8'had;
			8'h96: output_byte = 8'h35;
			8'h97: output_byte = 8'h85;
			8'h98: output_byte = 8'he2;
			8'h99: output_byte = 8'hf9;
			8'h9a: output_byte = 8'h37;
			8'h9b: output_byte = 8'he8;
			8'h9c: output_byte = 8'h1c;
			8'h9d: output_byte = 8'h75;
			8'h9e: output_byte = 8'hdf;
			8'h9f: output_byte = 8'h6e;
			8'ha0: output_byte = 8'h47;
			8'ha1: output_byte = 8'hf1;
			8'ha2: output_byte = 8'h1a;
			8'ha3: output_byte = 8'h71;
			8'ha4: output_byte = 8'h1d;
			8'ha5: output_byte = 8'h29;
			8'ha6: output_byte = 8'hc5;
			8'ha7: output_byte = 8'h89;
			8'ha8: output_byte = 8'h6f;
			8'ha9: output_byte = 8'hb7;
			8'haa: output_byte = 8'h62;
			8'hab: output_byte = 8'h0e;
			8'hac: output_byte = 8'haa;
			8'had: output_byte = 8'h18;
			8'hae: output_byte = 8'hbe;
			8'haf: output_byte = 8'h1b;
			8'hb0: output_byte = 8'hfc;
			8'hb1: output_byte = 8'h56;
			8'hb2: output_byte = 8'h3e;
			8'hb3: output_byte = 8'h4b;
			8'hb4: output_byte = 8'hc6;
			8'hb5: output_byte = 8'hd2;
			8'hb6: output_byte = 8'h79;
			8'hb7: output_byte = 8'h20;
			8'hb8: output_byte = 8'h9a;
			8'hb9: output_byte = 8'hdb;
			8'hba: output_byte = 8'hc0;
			8'hbb: output_byte = 8'hfe;
			8'hbc: output_byte = 8'h78;
			8'hbd: output_byte = 8'hcd;
			8'hbe: output_byte = 8'h5a;
			8'hbf: output_byte = 8'hf4;
			8'hc0: output_byte = 8'h1f;
			8'hc1: output_byte = 8'hdd;
			8'hc2: output_byte = 8'ha8;
			8'hc3: output_byte = 8'h33;
			8'hc4: output_byte = 8'h88;
			8'hc5: output_byte = 8'h07;
			8'hc6: output_byte = 8'hc7;
			8'hc7: output_byte = 8'h31;
			8'hc8: output_byte = 8'hb1;
			8'hc9: output_byte = 8'h12;
			8'hca: output_byte = 8'h10;
			8'hcb: output_byte = 8'h59;
			8'hcc: output_byte = 8'h27;
			8'hcd: output_byte = 8'h80;
			8'hce: output_byte = 8'hec;
			8'hcf: output_byte = 8'h5f;
			8'hd0: output_byte = 8'h60;
			8'hd1: output_byte = 8'h51;
			8'hd2: output_byte = 8'h7f;
			8'hd3: output_byte = 8'ha9;
			8'hd4: output_byte = 8'h19;
			8'hd5: output_byte = 8'hb5;
			8'hd6: output_byte = 8'h4a;
			8'hd7: output_byte = 8'h0d;
			8'hd8: output_byte = 8'h2d;
			8'hd9: output_byte = 8'he5;
			8'hda: output_byte = 8'h7a;
			8'hdb: output_byte = 8'h9f;
			8'hdc: output_byte = 8'h93;
			8'hdd: output_byte = 8'hc9;
			8'hde: output_byte = 8'h9c;
			8'hdf: output_byte = 8'hef;
			8'he0: output_byte = 8'ha0;
			8'he1: output_byte = 8'he0;
			8'he2: output_byte = 8'h3b;
			8'he3: output_byte = 8'h4d;
			8'he4: output_byte = 8'hae;
			8'he5: output_byte = 8'h2a;
			8'he6: output_byte = 8'hf5;
			8'he7: output_byte = 8'hb0;
			8'he8: output_byte = 8'hc8;
			8'he9: output_byte = 8'heb;
			8'hea: output_byte = 8'hbb;
			8'heb: output_byte = 8'h3c;
			8'hec: output_byte = 8'h83;
			8'hed: output_byte = 8'h53;
			8'hee: output_byte = 8'h99;
			8'hef: output_byte = 8'h61;
			8'hf0: output_byte = 8'h17;
			8'hf1: output_byte = 8'h2b;
			8'hf2: output_byte = 8'h04;
			8'hf3: output_byte = 8'h7e;
			8'hf4: output_byte = 8'hba;
			8'hf5: output_byte = 8'h77;
			8'hf6: output_byte = 8'hd6;
			8'hf7: output_byte = 8'h26;
			8'hf8: output_byte = 8'he1;
			8'hf9: output_byte = 8'h69;
			8'hfa: output_byte = 8'h14;
			8'hfb: output_byte = 8'h63;
			8'hfc: output_byte = 8'h55;
			8'hfd: output_byte = 8'h21;
			8'hfe: output_byte = 8'h0c;
			8'hff: output_byte = 8'h7d;
        endcase
    end

endmodule

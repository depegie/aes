`ifndef SCOREBOARD_SVH
`define SCOREBOARD_SVH

class scoreboard;

endclass

`endif

package tb_pkg;

    typedef struct {
        int         id;
        logic [7:0] data [$];
    } stream_t;

endpackage

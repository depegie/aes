`ifndef GENERATOR_SVH
`define GENERATOR_SVH

class generator;

endclass

`endif

`define AES256_CBC_ITER
`define S_AXIS_WIDTH 64
`define M_AXIS_WIDTH 64
`define S_AXIS_DELAY 0
`define M_AXIS_DELAY 0

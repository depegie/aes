package tb_pkg;

    typedef struct {
        int         id;
        logic [7:0] data [$];
    } packet_t;

endpackage

`define AES128_ECB_ITER_BEHAV
`define S_AXIS_WIDTH 64
`define M_AXIS_WIDTH 64
`define S_AXIS_DELAY 1
`define M_AXIS_DELAY 1

`include "aes_defines.svh"

module aes_inv_round_param #(
    parameter bit LAST = 0
)(
    input                          Enc,
    input  [`AES_BLOCK_SIZE-1 : 0] Input_block,
    output [`AES_BLOCK_SIZE-1 : 0] Output_block
);



endmodule

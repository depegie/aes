`ifndef MONITOR_SVH
`define MONITOR_SVH

class monitor;

endclass

`endif

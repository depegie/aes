`define AES_CBC_ITERATIVE
`define S_AXIS_DELAY 0
`define M_AXIS_DELAY 0

module aes_inv_sbox (
    input      [7 : 0] Input_byte,
    output reg [7 : 0] Output_byte
);
    always_comb begin
        case (Input_byte)
    		8'h00: Output_byte = 8'h52;
			8'h01: Output_byte = 8'h09;
			8'h02: Output_byte = 8'h6a;
			8'h03: Output_byte = 8'hd5;
			8'h04: Output_byte = 8'h30;
			8'h05: Output_byte = 8'h36;
			8'h06: Output_byte = 8'ha5;
			8'h07: Output_byte = 8'h38;
			8'h08: Output_byte = 8'hbf;
			8'h09: Output_byte = 8'h40;
			8'h0a: Output_byte = 8'ha3;
			8'h0b: Output_byte = 8'h9e;
			8'h0c: Output_byte = 8'h81;
			8'h0d: Output_byte = 8'hf3;
			8'h0e: Output_byte = 8'hd7;
			8'h0f: Output_byte = 8'hfb;
			8'h10: Output_byte = 8'h7c;
			8'h11: Output_byte = 8'he3;
			8'h12: Output_byte = 8'h39;
			8'h13: Output_byte = 8'h82;
			8'h14: Output_byte = 8'h9b;
			8'h15: Output_byte = 8'h2f;
			8'h16: Output_byte = 8'hff;
			8'h17: Output_byte = 8'h87;
			8'h18: Output_byte = 8'h34;
			8'h19: Output_byte = 8'h8e;
			8'h1a: Output_byte = 8'h43;
			8'h1b: Output_byte = 8'h44;
			8'h1c: Output_byte = 8'hc4;
			8'h1d: Output_byte = 8'hde;
			8'h1e: Output_byte = 8'he9;
			8'h1f: Output_byte = 8'hcb;
			8'h20: Output_byte = 8'h54;
			8'h21: Output_byte = 8'h7b;
			8'h22: Output_byte = 8'h94;
			8'h23: Output_byte = 8'h32;
			8'h24: Output_byte = 8'ha6;
			8'h25: Output_byte = 8'hc2;
			8'h26: Output_byte = 8'h23;
			8'h27: Output_byte = 8'h3d;
			8'h28: Output_byte = 8'hee;
			8'h29: Output_byte = 8'h4c;
			8'h2a: Output_byte = 8'h95;
			8'h2b: Output_byte = 8'h0b;
			8'h2c: Output_byte = 8'h42;
			8'h2d: Output_byte = 8'hfa;
			8'h2e: Output_byte = 8'hc3;
			8'h2f: Output_byte = 8'h4e;
			8'h30: Output_byte = 8'h08;
			8'h31: Output_byte = 8'h2e;
			8'h32: Output_byte = 8'ha1;
			8'h33: Output_byte = 8'h66;
			8'h34: Output_byte = 8'h28;
			8'h35: Output_byte = 8'hd9;
			8'h36: Output_byte = 8'h24;
			8'h37: Output_byte = 8'hb2;
			8'h38: Output_byte = 8'h76;
			8'h39: Output_byte = 8'h5b;
			8'h3a: Output_byte = 8'ha2;
			8'h3b: Output_byte = 8'h49;
			8'h3c: Output_byte = 8'h6d;
			8'h3d: Output_byte = 8'h8b;
			8'h3e: Output_byte = 8'hd1;
			8'h3f: Output_byte = 8'h25;
			8'h40: Output_byte = 8'h72;
			8'h41: Output_byte = 8'hf8;
			8'h42: Output_byte = 8'hf6;
			8'h43: Output_byte = 8'h64;
			8'h44: Output_byte = 8'h86;
			8'h45: Output_byte = 8'h68;
			8'h46: Output_byte = 8'h98;
			8'h47: Output_byte = 8'h16;
			8'h48: Output_byte = 8'hd4;
			8'h49: Output_byte = 8'ha4;
			8'h4a: Output_byte = 8'h5c;
			8'h4b: Output_byte = 8'hcc;
			8'h4c: Output_byte = 8'h5d;
			8'h4d: Output_byte = 8'h65;
			8'h4e: Output_byte = 8'hb6;
			8'h4f: Output_byte = 8'h92;
			8'h50: Output_byte = 8'h6c;
			8'h51: Output_byte = 8'h70;
			8'h52: Output_byte = 8'h48;
			8'h53: Output_byte = 8'h50;
			8'h54: Output_byte = 8'hfd;
			8'h55: Output_byte = 8'hed;
			8'h56: Output_byte = 8'hb9;
			8'h57: Output_byte = 8'hda;
			8'h58: Output_byte = 8'h5e;
			8'h59: Output_byte = 8'h15;
			8'h5a: Output_byte = 8'h46;
			8'h5b: Output_byte = 8'h57;
			8'h5c: Output_byte = 8'ha7;
			8'h5d: Output_byte = 8'h8d;
			8'h5e: Output_byte = 8'h9d;
			8'h5f: Output_byte = 8'h84;
			8'h60: Output_byte = 8'h90;
			8'h61: Output_byte = 8'hd8;
			8'h62: Output_byte = 8'hab;
			8'h63: Output_byte = 8'h00;
			8'h64: Output_byte = 8'h8c;
			8'h65: Output_byte = 8'hbc;
			8'h66: Output_byte = 8'hd3;
			8'h67: Output_byte = 8'h0a;
			8'h68: Output_byte = 8'hf7;
			8'h69: Output_byte = 8'he4;
			8'h6a: Output_byte = 8'h58;
			8'h6b: Output_byte = 8'h05;
			8'h6c: Output_byte = 8'hb8;
			8'h6d: Output_byte = 8'hb3;
			8'h6e: Output_byte = 8'h45;
			8'h6f: Output_byte = 8'h06;
			8'h70: Output_byte = 8'hd0;
			8'h71: Output_byte = 8'h2c;
			8'h72: Output_byte = 8'h1e;
			8'h73: Output_byte = 8'h8f;
			8'h74: Output_byte = 8'hca;
			8'h75: Output_byte = 8'h3f;
			8'h76: Output_byte = 8'h0f;
			8'h77: Output_byte = 8'h02;
			8'h78: Output_byte = 8'hc1;
			8'h79: Output_byte = 8'haf;
			8'h7a: Output_byte = 8'hbd;
			8'h7b: Output_byte = 8'h03;
			8'h7c: Output_byte = 8'h01;
			8'h7d: Output_byte = 8'h13;
			8'h7e: Output_byte = 8'h8a;
			8'h7f: Output_byte = 8'h6b;
			8'h80: Output_byte = 8'h3a;
			8'h81: Output_byte = 8'h91;
			8'h82: Output_byte = 8'h11;
			8'h83: Output_byte = 8'h41;
			8'h84: Output_byte = 8'h4f;
			8'h85: Output_byte = 8'h67;
			8'h86: Output_byte = 8'hdc;
			8'h87: Output_byte = 8'hea;
			8'h88: Output_byte = 8'h97;
			8'h89: Output_byte = 8'hf2;
			8'h8a: Output_byte = 8'hcf;
			8'h8b: Output_byte = 8'hce;
			8'h8c: Output_byte = 8'hf0;
			8'h8d: Output_byte = 8'hb4;
			8'h8e: Output_byte = 8'he6;
			8'h8f: Output_byte = 8'h73;
			8'h90: Output_byte = 8'h96;
			8'h91: Output_byte = 8'hac;
			8'h92: Output_byte = 8'h74;
			8'h93: Output_byte = 8'h22;
			8'h94: Output_byte = 8'he7;
			8'h95: Output_byte = 8'had;
			8'h96: Output_byte = 8'h35;
			8'h97: Output_byte = 8'h85;
			8'h98: Output_byte = 8'he2;
			8'h99: Output_byte = 8'hf9;
			8'h9a: Output_byte = 8'h37;
			8'h9b: Output_byte = 8'he8;
			8'h9c: Output_byte = 8'h1c;
			8'h9d: Output_byte = 8'h75;
			8'h9e: Output_byte = 8'hdf;
			8'h9f: Output_byte = 8'h6e;
			8'ha0: Output_byte = 8'h47;
			8'ha1: Output_byte = 8'hf1;
			8'ha2: Output_byte = 8'h1a;
			8'ha3: Output_byte = 8'h71;
			8'ha4: Output_byte = 8'h1d;
			8'ha5: Output_byte = 8'h29;
			8'ha6: Output_byte = 8'hc5;
			8'ha7: Output_byte = 8'h89;
			8'ha8: Output_byte = 8'h6f;
			8'ha9: Output_byte = 8'hb7;
			8'haa: Output_byte = 8'h62;
			8'hab: Output_byte = 8'h0e;
			8'hac: Output_byte = 8'haa;
			8'had: Output_byte = 8'h18;
			8'hae: Output_byte = 8'hbe;
			8'haf: Output_byte = 8'h1b;
			8'hb0: Output_byte = 8'hfc;
			8'hb1: Output_byte = 8'h56;
			8'hb2: Output_byte = 8'h3e;
			8'hb3: Output_byte = 8'h4b;
			8'hb4: Output_byte = 8'hc6;
			8'hb5: Output_byte = 8'hd2;
			8'hb6: Output_byte = 8'h79;
			8'hb7: Output_byte = 8'h20;
			8'hb8: Output_byte = 8'h9a;
			8'hb9: Output_byte = 8'hdb;
			8'hba: Output_byte = 8'hc0;
			8'hbb: Output_byte = 8'hfe;
			8'hbc: Output_byte = 8'h78;
			8'hbd: Output_byte = 8'hcd;
			8'hbe: Output_byte = 8'h5a;
			8'hbf: Output_byte = 8'hf4;
			8'hc0: Output_byte = 8'h1f;
			8'hc1: Output_byte = 8'hdd;
			8'hc2: Output_byte = 8'ha8;
			8'hc3: Output_byte = 8'h33;
			8'hc4: Output_byte = 8'h88;
			8'hc5: Output_byte = 8'h07;
			8'hc6: Output_byte = 8'hc7;
			8'hc7: Output_byte = 8'h31;
			8'hc8: Output_byte = 8'hb1;
			8'hc9: Output_byte = 8'h12;
			8'hca: Output_byte = 8'h10;
			8'hcb: Output_byte = 8'h59;
			8'hcc: Output_byte = 8'h27;
			8'hcd: Output_byte = 8'h80;
			8'hce: Output_byte = 8'hec;
			8'hcf: Output_byte = 8'h5f;
			8'hd0: Output_byte = 8'h60;
			8'hd1: Output_byte = 8'h51;
			8'hd2: Output_byte = 8'h7f;
			8'hd3: Output_byte = 8'ha9;
			8'hd4: Output_byte = 8'h19;
			8'hd5: Output_byte = 8'hb5;
			8'hd6: Output_byte = 8'h4a;
			8'hd7: Output_byte = 8'h0d;
			8'hd8: Output_byte = 8'h2d;
			8'hd9: Output_byte = 8'he5;
			8'hda: Output_byte = 8'h7a;
			8'hdb: Output_byte = 8'h9f;
			8'hdc: Output_byte = 8'h93;
			8'hdd: Output_byte = 8'hc9;
			8'hde: Output_byte = 8'h9c;
			8'hdf: Output_byte = 8'hef;
			8'he0: Output_byte = 8'ha0;
			8'he1: Output_byte = 8'he0;
			8'he2: Output_byte = 8'h3b;
			8'he3: Output_byte = 8'h4d;
			8'he4: Output_byte = 8'hae;
			8'he5: Output_byte = 8'h2a;
			8'he6: Output_byte = 8'hf5;
			8'he7: Output_byte = 8'hb0;
			8'he8: Output_byte = 8'hc8;
			8'he9: Output_byte = 8'heb;
			8'hea: Output_byte = 8'hbb;
			8'heb: Output_byte = 8'h3c;
			8'hec: Output_byte = 8'h83;
			8'hed: Output_byte = 8'h53;
			8'hee: Output_byte = 8'h99;
			8'hef: Output_byte = 8'h61;
			8'hf0: Output_byte = 8'h17;
			8'hf1: Output_byte = 8'h2b;
			8'hf2: Output_byte = 8'h04;
			8'hf3: Output_byte = 8'h7e;
			8'hf4: Output_byte = 8'hba;
			8'hf5: Output_byte = 8'h77;
			8'hf6: Output_byte = 8'hd6;
			8'hf7: Output_byte = 8'h26;
			8'hf8: Output_byte = 8'he1;
			8'hf9: Output_byte = 8'h69;
			8'hfa: Output_byte = 8'h14;
			8'hfb: Output_byte = 8'h63;
			8'hfc: Output_byte = 8'h55;
			8'hfd: Output_byte = 8'h21;
			8'hfe: Output_byte = 8'h0c;
			8'hff: Output_byte = 8'h7d;
        endcase
    end

endmodule

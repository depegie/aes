`ifndef DRIVER_SVH
`define DRIVER_SVH

class driver;

endclass

`endif
